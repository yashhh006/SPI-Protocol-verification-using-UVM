typedef uvm_sequencer #(apb_tx) spi_sqr;